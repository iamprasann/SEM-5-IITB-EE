Prasann Viswanathan 190070047 RC Low-pass Filter

r1 1 2 10k
c1 2 0 0.1u
v_in 1 0 dc 0 ac 1

*analysis command
.ac dec 10 1 10k
.control
run

*display commands
plot vdb(2)
.endc
.end 