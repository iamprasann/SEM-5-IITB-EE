Prasann Viswanathan 190070047 RC Integrator

r1 1 2 10k
c1 2 0 0.1u
*v_in 1 0 pulse(0 5 0.1u 0 0 10m 20m)
v_in 1 0 pulse(0 5 0.1u 0 0 1m 2m)

*analysis command
*.tran 10u 40m
.tran 10u 10m
.control
run

*display commands
plot v(2) v(1)
.endc
.end 