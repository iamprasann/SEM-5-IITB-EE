Prasann Viswanathan 190070047 NMOS Common Source Amp Experiment

.model mos_model nmos Level=1 Vto=1 KP=100u w=10u L=1u
+ Gamma=0 Phi=0.65 Lambda=0.0

vin 3 0 sin(0 50m 1k 0 0)
vdd 1 0 12
v_t 1 2 0
r1 1 g 8.2k
r2 g 0 3.3k
rd 2 d 3.3k
rs s 0 1k
m1 d g s 0 mos_model
c1 g 3 10u
c2 s 0 100u

*analysis commands
.tran 10u 20ms
.control
run

*display commands
plot v(3)
plot v(d)
.endc 
.end