Prasann Viswanathan 190070047 NMOS Current Mirror Current Source

.model mos_model nmos Level=1 Vto=1 KP=100u w=10u L=1u
+ Gamma=0 Phi=0.65 Lambda=0.0

vdd 1 0 12
m1 2 2 0 0 mos_model
m2 3 2 0 0 mos_model
v0 3 0 0
r 1 2 8.2k

*analysis commands
.dc v0 1 5 0.2
.control
run

*display commands
plot -i(v0)
plot -i(vdd)
print -i(v0)
print -i(vdd)
.endc
.end