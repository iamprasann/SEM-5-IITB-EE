Prasann Viswanathan 190070047 regulated BJT series

.include zener_B.txt

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

.model SL100 NPN IS=100f BF=80 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=100 RE=1 RC=10
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

v_in 1 0
q1 3 4 5 bc547a
q2 1 3 2 SL100
rc 1 3 1k
r1 2 4 10.2k
r2 4 0 14.8k
rl 2 0 1k
x1 0 5 DI_1N4734A

*analysis command
.dc Vin 15 25 0.5

.control
run

*display commands
print v(1) v(2) v(3) v(4) v(5)
plot v(1) v(2) v(3) v(4) v(5)

.endc
.end