Prasann Viswanathan 190070047 NMOS Characteristics

.model NXYAA5U nmos Level=1 Vto=0.7 KP=80u w=10u L=1u
+ Gamma=0 Phi=0.65 Lambda=0.0

vgs 2 0 0
v2 1 0 0
rd 1 3 2.2k
m1 3 2 0 0 NXYAA5U

*analysis commands
.dc v2 0 50 0.02 Vgs 2 5 1
.control
run

*display commands
plot -i(v2)
.endc
.end