Prasann Viswanathan 190070047 BJT Current Source

.include zener_B.txt
.model bc557a PNP IS=10f BF=100 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

q1 4 3 2 bc557a
vcc 1 0 12
vl 5 0 0
xz 3 1 DI_1N4734A
re 1 2 4.7k
rb 3 0 2.2k
rl 4 5 1k

*analysis commands
.op 
.control
run

*display commands
print i(vl) v(2) v(3) v(4)
.endc
.end