Prasann Viswanathan 190070047 Common Emitter

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

q1 c b e bc547a
vc 3 c 0
vb 2 b 0
ve e 1 0
vcc 4 0 12
re 1 0 1k
rc 4 3 1.2k
r1 4 2 10k
r2 2 0 2.2k

*analysis commands
.op
.control
run

*display commands
print i(vb) i(vc) v(b) v(c) v(e)
.endc
.end