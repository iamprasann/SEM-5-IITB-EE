Prasann Viswanathan 190070047 BJT Current Mirror

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

q1 2 2 0 bc547a
q2 3 2 0 bc547a
vcc 1 0 12
vo 3 0 1
r 1 2 10k

*analysis commands
.op
.control
run 

*display commands
print i(vcc) i(vo) v(2)
.endc
.end